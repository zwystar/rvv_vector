module vec_dec
    #(
        parameter XLEN = 512,
        parameter SEW  = 32
    )
    (
    input  clk,    // Clock
    input  clk_en, // Clock Enable
    input  rst_n,  // Asynchronous reset active low
    
    input 
);



endmodule
